module maindec (
        input  wire [5:0] opcode,
        output wire       branch,
        output wire       jump,
        output wire       jal,
        output wire       reg_dst,
        output wire       we_reg,
        output wire       alu_src,
        output wire       we_dm,
        output wire       dm2reg,
        output wire [1:0] alu_op,
        output wire       iack,
        output wire       rfe
    );

    reg [11:0] ctrl;

    assign {branch, jump, reg_dst, we_reg, alu_src, we_dm, dm2reg, alu_op, jal, iack, rfe} = ctrl;

    always @ (opcode) begin
        case (opcode)
            6'b00_0000: ctrl = 12'b0_0_1_1_0_0_0_10_0_0_0; // R-type
            6'b00_1000: ctrl = 12'b0_0_0_1_1_0_0_00_0_0_0; // ADDI
            6'b00_0100: ctrl = 12'b1_0_0_0_0_0_0_01_0_0_0; // BEQ
            6'b00_0010: ctrl = 12'b0_1_0_0_0_0_0_00_0_0_0; // J
            6'b00_0011: ctrl = 12'b0_1_0_1_0_0_0_00_1_0_0; // JAL
            6'b10_1011: ctrl = 12'b0_0_0_0_1_1_0_00_0_0_0; // SW
            6'b10_0011: ctrl = 12'b0_0_0_1_1_0_1_00_0_0_0; // LW
            6'b11_0000: ctrl = 12'b0_0_0_0_0_0_0_00_0_1_0; // IACK
            6'b11_0001: ctrl = 12'b0_0_0_0_0_0_0_00_0_1_1; // RFE
            default:    ctrl = 12'bx_x_x_x_x_x_x_xx_x_x_x;
        endcase
    end

endmodule
